`default_nettype none
module top (input wire clk);
    reg test = 0;
endmodule
